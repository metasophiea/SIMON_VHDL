library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.textio.all; 
use work.printerlib.all;

entity messageEncrypter is
    port(
        instance: in std_logic_vector(7 downto 0);
        method: in std_logic_vector(3 downto 0);
        keyIn: in std_logic_vector(255 downto 0);
        messageIn: in std_logic_vector(127 downto 0);
        messageOut: out std_logic_vector(127 downto 0)
    );
end messageEncrypter;

architecture behaviour of messageEncrypter is
-- //////// //////// //////// //////// //////// //////// //////// ////////
     -- tools
    function morph_Z(Z: std_logic_vector)
    return std_logic_vector is variable Z_manipulator: std_logic_vector(61 downto 0) := Z;
    begin return Z_manipulator(Z_manipulator'length-2 downto 0) & Z_manipulator(Z_manipulator'length-1);
    end function;

    function rightRotate(logic: std_logic_vector; amount: integer)
    return std_logic_vector is  variable temp: std_logic_vector(logic'length-1 downto 0) := logic;
    begin
        for a in 0 to amount-1 loop  temp := temp(0) & temp(temp'length-1 downto 1);  end loop;
        return temp;
    end function;

    function leftRotate(logic: std_logic_vector; amount: integer)
    return std_logic_vector is  variable temp: std_logic_vector(logic'length-1 downto 0) := logic;
    begin
        for a in 0 to amount-1 loop  temp := temp(temp'length-2 downto 0) & temp(temp'length-1); end loop;
        return temp;
    end function;
    
    -- main encryptor work function
    function encryptor_workFunction(messageIn, keyIn: std_logic_vector; segmentLength, keyLength, keySegments: integer)
    return std_logic_vector is
        variable combiner: std_logic_vector(127 downto 0) := (others => '0');
        variable x, y, holder, temp, key: std_logic_vector(63 downto 0) := (others => '0');
    begin
        -- aquire parts
        x(segmentLength-1 downto 0) := messageIn((2*segmentLength)-1 downto segmentLength);
        y(segmentLength-1 downto 0) := messageIn(segmentLength-1 downto 0);
        key(segmentLength-1 downto 0) := keyIn(keyLength-1-(segmentLength*(keySegments-1)) downto keyLength-segmentLength-(segmentLength*(keySegments-1)));
    
        -- encryption
        holder := x;
        temp(segmentLength-1 downto 0) := leftRotate(x(segmentLength-1 downto 0),1) and leftRotate(x(segmentLength-1 downto 0),8);
        temp(segmentLength-1 downto 0) := temp(segmentLength-1 downto 0) xor y(segmentLength-1 downto 0);
        temp(segmentLength-1 downto 0) := temp(segmentLength-1 downto 0) xor leftRotate(x(segmentLength-1 downto 0),2);
        temp(segmentLength-1 downto 0) := temp(segmentLength-1 downto 0) xor key(segmentLength-1 downto 0);
        x := temp; y := holder;
    
        -- recombination
        combiner((2*segmentLength)-1 downto segmentLength) := x(segmentLength-1 downto 0);
        combiner(segmentLength-1 downto 0) := y(segmentLength-1 downto 0); 
        return combiner;
    end function; 

    -- main encryptor
    function encrypt(messageIn, keyIn, method: std_logic_vector)
    return std_logic_vector is
        variable segmentLength, keyLength, keySegments: integer := 0;
    begin
        case (std_logic_vector(method)) is
            when "0000" => segmentLength := 16; keySegments := 4; keyLength := 64; 
            when "0001" => segmentLength := 24; keySegments := 3; keyLength := 72; 
            when "0010" => segmentLength := 24; keySegments := 4; keyLength := 96; 
            when "0011" => segmentLength := 32; keySegments := 3; keyLength := 96; 
            when "0100" => segmentLength := 32; keySegments := 4; keyLength := 128;
            when "0101" => segmentLength := 48; keySegments := 2; keyLength := 96; 
            when "0110" => segmentLength := 48; keySegments := 3; keyLength := 144;
            when "0111" => segmentLength := 64; keySegments := 2; keyLength := 128;
            when "1000" => segmentLength := 64; keySegments := 3; keyLength := 192;
            when "1001" => segmentLength := 64; keySegments := 4; keyLength := 256;
            when others => segmentLength := 64; keySegments := 4; keyLength := 256;
        end case; 
		
		return encryptor_workFunction(messageIn, keyIn, segmentLength, keyLength, keySegments);
    end function;

begin
-- //////// //////// //////// //////// //////// //////// //////// ////////
    process(messageIn, keyIn, method) 
    begin 
        case method is
            when "0000" => if to_integer(unsigned(instance)) > (32-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "0001" => if to_integer(unsigned(instance)) > (36-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "0010" => if to_integer(unsigned(instance)) > (36-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "0011" => if to_integer(unsigned(instance)) > (42-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "0100" => if to_integer(unsigned(instance)) > (44-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "0101" => if to_integer(unsigned(instance)) > (52-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "0110" => if to_integer(unsigned(instance)) > (54-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "0111" => if to_integer(unsigned(instance)) > (68-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "1000" => if to_integer(unsigned(instance)) > (69-1) then messageOut <= messageIn; else messageOut <= encrypt(messageIn,keyIn,method); end if;
            when "1001" => messageOut <= encrypt(messageIn,keyIn,method);
            when others =>  messageOut <= messageIn;
        end case;
    end process;
end behaviour;