library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.textio.all; 
use work.printerlib.all;

-- Methods | messageLength/keyLength | keySegmentLength | keySegments | messageSegments | messageSegmentLength | cryptLoopCount | Zselect
-- 0000    | 32/64                   | 16               | 4           | 2               | 16                   | 32             | 0

entity simon is
    port(
        mode: in std_logic;
        keyIn: in std_logic_vector(63 downto 0) := (others => '0');
        messageIn: in std_logic_vector(31 downto 0);
        messageOut: out std_logic_vector(31 downto 0) := (others => '0')
    );
end simon;

architecture behaviour of simon is
-- //////// //////// //////// //////// //////// //////// //////// ////////
    -- declare constants
    constant maxCryptLoopCount : integer := 32;

    -- declare components
    component keyExpander
        port(
            Z: in std_logic_vector(61 downto 0);
            keyIn: in std_logic_vector(63 downto 0);
            keyOut: out std_logic_vector(63 downto 0);
            returnZ: out std_logic_vector(61 downto 0)
        );
    end component;

    component messageEncrypter is
        port(
            keyIn: in std_logic_vector(63 downto 0);
            messageIn: in std_logic_vector(31 downto 0);
            messageOut: out std_logic_vector(31 downto 0)
        );
    end component;

    component messageDecrypter is
        port(
            keyIn: in std_logic_vector(63 downto 0);
            messageIn: in std_logic_vector(31 downto 0);
            messageOut: out std_logic_vector(31 downto 0)
        );
    end component;  

    -- declare Z's
    signal Z_0: std_logic_vector(61 downto 0) := "11111010001001010110000111001101111101000100101011000011100110";

    -- internal signals
    type morphingZ_type is array (0 to (maxCryptLoopCount-1)) of std_logic_vector(61 downto 0);
    signal morphingZ: morphingZ_type := ( others => std_logic_vector(to_unsigned(0,62)) );

    type morphingKey_type is array (0 to (maxCryptLoopCount-1)) of std_logic_vector(63 downto 0);
    signal morphingKey: morphingKey_type := ( others => std_logic_vector(to_unsigned(0,64)) );

    type morphingMessage_type is array (0 to maxCryptLoopCount) of std_logic_vector(31 downto 0); 
    signal morphingEncryptMessage: morphingMessage_type := ( others => std_logic_vector(to_unsigned(0,32)) );
    signal morphingDecryptMessage: morphingMessage_type := ( others => std_logic_vector(to_unsigned(0,32)) );

begin
    -- connect inputs
    morphingKey(0) <= keyIn;
    morphingEncryptMessage(0) <= messageIn;
    morphingDecryptMessage(0) <= messageIn;

    -- select Z baised on selected method
    morphingZ(0) <= Z_0;

-- generate and connect components
    keyExpansion_generation:for a in 0 to (maxCryptLoopCount-2) generate
        keyExpansion: keyExpander port map(    
            Z => morphingZ(a),
            returnZ => morphingZ(a+1),
            keyIn => morphingKey(a),
            keyOut => morphingKey(a+1)
        ); 
    end generate; 

    encrypterDecrypter_generation:for a in 0 to (maxCryptLoopCount-1) generate
        encryptMessage: messageEncrypter port map(
            keyIn => morphingKey(a),
            messageIn => morphingEncryptMessage(a),
            messageOut => morphingEncryptMessage(a+1)
        );

        decryptMessage: messageDecrypter port map(
            keyIn => morphingKey((maxCryptLoopCount-1)-a),
            messageIn => morphingDecryptMessage(a),
            messageOut => morphingDecryptMessage(a+1)
        );
    end generate;

    -- connect output
    messageOut <= morphingEncryptMessage(maxCryptLoopCount) when mode = '0' else morphingDecryptMessage(maxCryptLoopCount);
end behaviour;